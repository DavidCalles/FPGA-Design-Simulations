library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

package common is    -- untested...

    type regArray_t is array (1 to 7) of unsigned(15 downto 0);
 
 end common;
 
 package body common is

 end common;