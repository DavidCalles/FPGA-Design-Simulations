/* cpu.v:
 *
 * CPU implementation
 * 
 */

module CPU(/*AUTOARG*/
   // Outputs
   DATA_O, ADDR, RD, WR,
   // Inputs
   DATA_I, CLK, RST
   );
   input [15:0]  DATA_I;
   output [15:0] DATA_O;
   output [15:0] ADDR;
   output 	 RD;
   output 	 WR;
   
   input 	 CLK;
   input 	 RST;
 
   reg [15:0] 	 IR;
   reg [15:0] 	 MAR;
   reg [10:0] 	 CAR,CAR_next;
   wire [10:0] 	 EXT_ADRS;
   
   wire [15:0] 	 ABUS,BBUS,FOUT;
   wire 	 LDMAR,LDIR,RFMUX,DMUX;
	    
   wire [10:0] MUX1_OUT;
   wire MUX2_OUT;

   /* Status flag registers, and wires */
   reg 		 Z,S,C,V;
   wire 	 ZOUT,SOUT,COUT,VOUT;
   wire          UPZ,UPS,UPC,UPV;
 	 
   
   /* Buffer address register, and data out signals */
   assign ADDR = MAR;
   assign DATA_O = FOUT;
   

   /* Instantiate microcode ROM */
   wire [43:0]  ROM_out;

   MICROCODE_ROM MICROCODE_ROM1(
      .ADDR_in(CAR),
      .ROM_out(ROM_out));

   wire [ 2:0]  ASEL;
   wire [ 2:0]  BSEL;
   wire [ 2:0]  DSEL;
   wire [ 3:0]  FSEL;
   wire [ 3:0]  UPDF;
   wire         MUX1;
   wire [ 3:0]  MUX2;
   wire [15:0]  DATA;
   wire [ 5:0]  MISC;

   assign                 ASEL = ROM_out[43:41];    // bit size:3
   assign                 BSEL = ROM_out[40:38];    // bit size:3
   assign                 DSEL = ROM_out[37:35];    // bit size:3
   assign                 FSEL = ROM_out[34:31];    // bit size:4
   assign                 UPDF = ROM_out[30:27];    // bit size:4
   assign                 MUX1 = ROM_out[26];       // bit size:1
   assign                 MUX2 = ROM_out[25:22];    // bit size:4
   assign                 DATA = ROM_out[21: 6];    // bit size:16
   assign                 MISC = ROM_out[ 5: 0];    // bit size:6

   /* Split out the MISC field */
   assign RD    = MISC[0];
   assign WR    = MISC[1];
   assign LDMAR = MISC[2];
   assign LDIR  = MISC[3];
   assign RFMUX = MISC[4];
   assign DMUX  = MISC[5];

   /* Split out Update Flags field */
   assign UPZ   = UPDF[3];
   assign UPS   = UPDF[2];
   assign UPC   = UPDF[1];
   assign UPV   = UPDF[0];
   
   /* Instantiate Register file */
   REGFILE REGFILE1(   // Outputs
		       .ABUS(ABUS),
		       .BBUS(BBUS),
		       // Inputs
		       .ASEL(RFMUX ? IR[8:6] : ASEL),
		       .BSEL(RFMUX ? IR[5:3] : BSEL),
		       .DSEL(RFMUX ? IR[2:0] : DSEL),
		       .DIN(DMUX ? DATA    : DATA_I),
		       .RIN(FOUT),
		       .CLK(CLK),
		       .RST(RST));
      
   /* Instantiate ALU */
   ALU ALU1(// Outputs
	    .FOUT(FOUT),
	    .C(COUT), .Z(ZOUT), .S(SOUT), .V(VOUT),
	    // Inputs
	    .ABUS(ABUS),
	    .BBUS(BBUS),
	    .FSEL(FSEL),
	    .CIN(C));

   /* ALU Flag updating */
   always @(posedge CLK or negedge RST)
     if(RST==1'b0) begin
	Z   <= 0;
	S   <= 0;
	C   <= 0;
	V   <= 0;
	MAR <= 0;
	IR  <= 0;
     end else begin
	if(UPZ) begin
	   Z <= ZOUT;
	end

	if(UPS) begin
	   S <= SOUT;
	end
	
	if(UPC) begin
	   C <= COUT;
	end
	
	if(UPV) begin
	   V <= VOUT;
	end

	if(LDMAR) begin
	   MAR <= ABUS;
	end

	if(LDIR) begin
	   IR <= DATA_I;
	end
     end

   /* Sequencer logic -- Implement your logic for CAR generation here */

   /* Muxes */
   assign EXT_ADRS = {1'b0, IR[15:9], 3'b000};

   always @ (posedge CLK or negedge RST or MUX2_OUT or MUX1_OUT)
   begin
      if (RST == 1'b0)
         CAR <= 0;
      else begin
         if(MUX2_OUT == 1'b0) 
            CAR <= CAR+1;  
         else if(MUX2_OUT) 
            CAR <= MUX1_OUT; 
      end 
   end   

assign MUX1_OUT = MUX1 == 1'b0 ? DATA[10:0] :
                  MUX1 == 1'b1 ? DATA_I[10:0] : 1'b0;

assign MUX2_OUT = MUX2 == 4'b0000 ? 1'b0 :
                  MUX2 == 4'b0001 ? 1'b1 :
                  MUX2 == 4'b0010 ? C : 
                  MUX2 == 4'b0011 ? ~C :
                  MUX2 == 4'b0100 ? Z :
                  MUX2 == 4'b0101 ? ~Z :
                  MUX2 == 4'b0110 ? S :
                  MUX2 == 4'b0111 ? ~S :
                  MUX2 == 4'b1000 ? V :
                  MUX2 == 4'b1001 ? ~V :
                  MUX2 == 4'b1010 ? S ^ V :
                  MUX2 == 4'b1011 ? ~(S^V) : 1'b0;
   
endmodule
	 
