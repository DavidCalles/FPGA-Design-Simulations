-- ALU entity